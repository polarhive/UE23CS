module NOT(input a, output y);
    assign y = !a;
endmodule