module main;
  initial 
    begin
      $display("Hello World");
      $finish ;
    end
endmodule
